`timescale 1ns / 1ps

module memory #(
    parameter MEMORY_SIZE = 262143
) (
    input clk,
    input we,
    input [31:0] addr,
    output logic [31:0] r_data,
    input [31:0] w_data);
    
(* ram_style = "block" *) logic [31:0] mem [0:MEMORY_SIZE];
    
    //initial $readmemb("read.coe", mem);
    
    initial begin
        mem[0] = 32'b01000011000000000000000000000000;
        mem[1] = 32'b00111111011001100110011001100110;
        mem[2] = 32'b00111110010011001100110011001101;
        mem[3] = 32'b01000011000101100000000000000000;
        mem[4] = 32'b11000011000101100000000000000000;
        mem[5] = 32'b00111101110011001100110011001101;
        mem[6] = 32'b11000000000000000000000000000000;
        mem[7] = 32'b00111011100000000000000000000000;
        mem[8] = 32'b01000001101000000000000000000000;
        mem[9] = 32'b00111101010011001100110011001101;
        mem[10] = 32'b00111110100000000000000000000000;
        mem[11] = 32'b01000001001000000000000000000000;
        mem[12] = 32'b00111110100110011001100110011010;
        mem[13] = 32'b01000011011111110000000000000000;
        mem[14] = 32'b00111111000000000000000000000000;
        mem[15] = 32'b00111110000110011001100110011010;
        mem[16] = 32'b01000000010010010000111111011011;
        mem[17] = 32'b01000001111100000000000000000000;
        mem[18] = 32'b01000001011100000000000000000000;
        mem[19] = 32'b00111000110100011011011100010111;
        mem[20] = 32'b01001100101111101011110000100000;
        mem[21] = 32'b01001110011011100110101100101000;
        mem[22] = 32'b10111101110011001100110011001101;
        mem[23] = 32'b00111100001000111101011100001010;
        mem[24] = 32'b10111110010011001100110011001101;
        mem[25] = 32'b01000000000000000000000000000000;
        mem[26] = 32'b11000011010010000000000000000000;
        mem[27] = 32'b01000011010010000000000000000000;
        mem[28] = 32'b00111100100011101111101000110101;
        mem[29] = 32'b10111111100000000000000000000000;
        mem[30] = 32'b00111111100000000000000000000000;
        mem[31] = 32'b00000000000000000000000000000000;
        mem[32] = 32'b00000000000000000000000000000000;
        mem[33] = 32'b00111111100000000000000000000000;
        mem[34] = 32'b01000000000000000000000000000000;
        mem[35] = 32'b01001011000000000000000000000000;
        mem[36] = 32'b01000001001000000000000000000000;
        mem[37] = 32'b00111111010010010000111111011011;
        mem[38] = 32'b00111111110010010000111111011011;
        mem[39] = 32'b01000000010010010000111111011011;
        mem[40] = 32'b01000000110010010000111111011011;
        mem[41] = 32'b00111110001010101010101010101100;
        mem[42] = 32'b00111100000010001000011001100110;
        mem[43] = 32'b00111001010011010110010010110110;
        mem[44] = 32'b00111111000000000000000000000000;
        mem[45] = 32'b00111101001010101010011110001001;
        mem[46] = 32'b00111010101100111000000100000110;
        mem[47] = 32'b00111110111000000000000000000000;
        mem[48] = 32'b01000000000111000000000000000000;
        mem[49] = 32'b00111110101010101010101010101010;
        mem[50] = 32'b00111110010011001100110011001101;
        mem[51] = 32'b00111110000100100100100100100101;
        mem[52] = 32'b00111101111000111000111000111000;
        mem[53] = 32'b00111101101101111101011001101110;
        mem[54] = 32'b00111101011101011110011111000101;
        mem[55] = 32'b00000000000000000000000000000000;
        mem[56] = 32'b00000000000000000000000000000000;
        mem[57] = 32'b00000000000000000000000000000000;
        mem[58] = 32'b00000000000000000000000000000000;
        mem[59] = 32'b00000000000000000000000000000000;
        mem[60] = 32'b00000000000000000000000000000000;
        mem[61] = 32'b00000000000000000000000000000000;
        mem[62] = 32'b00000000000000000000000000000000;
        mem[63] = 32'b00000000000000000000000000000000;
        mem[64] = 32'b00000000000000000000000000000000;
        mem[65] = 32'b00000000000000000000000000000000;
        mem[66] = 32'b00000000000000000000000000000000;
        mem[67] = 32'b00000000000000000000000000000000;
        mem[68] = 32'b00000000000000000000000000000000;
        mem[69] = 32'b00000000000000000000000000000000;
        mem[70] = 32'b00000000000000000000000000000000;
        mem[71] = 32'b00000000000000000000000000000000;
        mem[72] = 32'b00000000000000000000000000000000;
        mem[73] = 32'b00000000000000000000000000000000;
        mem[74] = 32'b00000000000000000000000000000000;
        mem[75] = 32'b00000000000000000000000000000000;
        mem[76] = 32'b00000000000000000000000000000000;
        mem[77] = 32'b00000000000000000000000000000000;
        mem[78] = 32'b00000000000000000000000000000000;
        mem[79] = 32'b00000000000000000000000000000000;
        mem[80] = 32'b00000000000000000000000000000000;
        mem[81] = 32'b00000000000000000000000000000000;
        mem[82] = 32'b00000000000000000000000000000000;
        mem[83] = 32'b00000000000000000000000000000000;
        mem[84] = 32'b00000000000000000000000000000000;
        mem[85] = 32'b00000000000000000000000000000000;
        mem[86] = 32'b00000000000000000000000000000000;
        mem[87] = 32'b00000000000000000000000000000000;
        mem[88] = 32'b00000000000000000000000000000000;
        mem[89] = 32'b00000000000000000000000000000000;
        mem[90] = 32'b00000000000000000000000000000000;
        mem[91] = 32'b00000000000000000000000000000000;
        mem[92] = 32'b00000000000000000000000000000000;
        mem[93] = 32'b00000000000000000000000000000000;
        mem[94] = 32'b00000000000000000000000000000000;
        mem[95] = 32'b00000000000000000000000000000000;
        mem[96] = 32'b00000000000000000000000000000000;
        mem[97] = 32'b00000000000000000000000000000000;
        mem[98] = 32'b00000000000000000000000000000000;
        mem[99] = 32'b00000000000000000000000000000000;
    end
    
    always @(posedge clk) begin
        if (we) mem[addr] <= w_data;
        r_data <= mem[addr];
    end
endmodule
